-- Boost Software License - Version 1.0 - August 17th, 2003 Timo Sarkar, Igel
--
-- Permission is hereby granted, free of charge, to any person or organization
-- obtaining a copy of the software and accompanying documentation covered by
-- this license (the "Software") to use, reproduce, display, distribute,
-- execute, and transmit the Software, and to prepare derivative works of the
-- Software, and to permit third-parties to whom the Software is furnished to
-- do so, all subject to the following:
--
-- The copyright notices in the Software and this entire statement, including
-- the above license grant, this restriction and the following disclaimer,
-- must be included in all copies of the Software, in whole or in part, and
-- all derivative works of the Software, unless such copies or derivative
-- works are solely in the form of machine-executable object code generated by
-- a source language processor.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE, TITLE AND NON-INFRINGEMENT. IN NO EVENT
-- SHALL THE COPYRIGHT HOLDERS OR ANYONE DISTRIBUTING THE SOFTWARE BE LIABLE
-- FOR ANY DAMAGES OR OTHER LIABILITY, WHETHER IN CONTRACT, TORT OR OTHERWISE,
-- ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
-- DEALINGS IN THE SOFTWARE.

library STD;
use STD.textio.all;

package pkg_readline is
    procedure igel_printline( li: string );
    procedure igel_readline( prompt: string: eof_detected: out boolean; l: inout line );
end package pkg_readline;

package body pkg_readline is 
    type charfile is file of character;
    file stdout_char: charfile open write_mode is "STD_OUTPUT";

    procedure igel_printstr( l: string ) is 
    begin
        for i in l'range loop
            write( stdout_char, l( i ) );
        end loop;
    end procedure igel_printstr;
    
    procedure igel_printline( l: string ) is
    begin
        igel_printstr( l );
        write( stdout_char, LF );
    end procedure igel_printline;

    procedure igel_readline( prompt: string; eof_detected: out boolean; l: inout line ) is 
    begin
        igel_printstr( prompt );
        if endfile( input ) then
            eof_detected := true;
        else
            readline( input, 1 );
            eof_detected := false;
        end if;
    end procedure igel_readline;
end package body pkg_readline; 
