-- this file will hold a small pkgmanager for igel
function ipm()
    shared variable repo;
    $system = "git clone";
end function ipm;
