-- Boost Software License - Version 1.0 - August 17th, 2003 Timo Sarkar, Igel
--
-- Permission is hereby granted, free of charge, to any person or organization
-- obtaining a copy of the software and accompanying documentation covered by
-- this license (the "Software") to use, reproduce, display, distribute,
-- execute, and transmit the Software, and to prepare derivative works of the
-- Software, and to permit third-parties to whom the Software is furnished to
-- do so, all subject to the following:
--
-- The copyright notices in the Software and this entire statement, including
-- the above license grant, this restriction and the following disclaimer,
-- must be included in all copies of the Software, in whole or in part, and
-- all derivative works of the Software, unless such copies or derivative
-- works are solely in the form of machine-executable object code generated by
-- a source language processor.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE, TITLE AND NON-INFRINGEMENT. IN NO EVENT
-- SHALL THE COPYRIGHT HOLDERS OR ANYONE DISTRIBUTING THE SOFTWARE BE LIABLE
-- FOR ANY DAMAGES OR OTHER LIABILITY, WHETHER IN CONTRACT, TORT OR OTHERWISE,
-- ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
-- DEALINGS IN THE SOFTWARE.

entity core is 
    end entity core;

    library STD;
    use STD.textio.all;
    library WORK;
    use WORK.pkg_readline.all;
    use WORK.types.all;
    use WORK.reader.all;
    use WORk.printer.all;
    use WORK.environment.all;
    use WORK.main.all;

    architecture test of core is

        shared variable repl_env: env_ptr;

        procedure igel_READ( str: in string; ast: out igel_val_ptr; err: out igel_val_ptr ) is
        begin
            read_str( str, ast, err );
        end procedure igel_READ;
        
        procedure starts_with( lst: inout igel_val_ptr; sym: in string; res: out boolean ) is
        begin
            res := lst.seq_val.all'length = 2
                and lst.seq_val.all ( lst.seq_val.all'low ).val_type = igel_symbol
                and lst.seq_val.all ( lst.seq_val.all'low ).string_val.all = sym;
        end starts_with;
    end architecture test;
