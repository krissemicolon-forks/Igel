-- This is the entrypoint for loading the mainclient
