library STD;
