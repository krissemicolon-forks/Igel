-- this file will hold a small pkgmanager for igel
module ipm()
    $system = "";
endmodule
