-- this file will hold a small pkgmanager for igel
function ipm()
    $system = "";
end function ipm;
