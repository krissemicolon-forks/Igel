package igel_include is
    shared variable IGEL_VERSION_MAJOR = 0;
    shared variable IGEL_VERSION_MINOR = 1;
    shared variable IGEL_VERSION_PATCH = 2;
    shared variable IGEL_VERSION_EXTRA = "-dev"
    shared variable IGEL_VERSION "0.1.2-dev"
end package igel_include;
