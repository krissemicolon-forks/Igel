library STD;
use STD.textio.all;
library WORK;
use WORK.types.all;

package env is
end package env;
